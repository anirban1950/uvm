package agt_pkg;
   import uvm_pkg::*;
  `include "packet.sv"
  `include "packet2.sv"
  `include "monitor.sv"
  `include "driver.sv"
  `include "agent.sv"
endpackage
