package test_pkg;
   import uvm_pkg::*;
   import agt_pkg::*;
  `include "base_seq.sv"
  `include "env.sv"
  `include "test_base.sv"
  `include "test1.sv"
  `include "test2.sv"
endpackage
