// Code your testbench here
// or browse Examples
`include "agt_pkg.sv"
`include "test_pkg.sv"
`include "top.sv"